`timescale 1ns/1ps

module test_alu;
reg[31:0] instruction;
reg[31:0] regA;
reg[31:0] regB;
wire[2:0] flags;
wire[31:0] result;
alu dut(.instruction(instruction), .regA(regA), .regB(regB), .flags(flags), .result(result));
initial begin

    #10
    $display("add");
    instruction = 32'b000000_00001_00000_00000_00000_100000;
    regA = 32'h00000001;
    regB = 32'h00000003; //3+1
    $monitor("instruction: %b\nregA: %b\nregB: %b\nflags: %b\nresult: %b\n", 
            instruction, regA, regB, flags, result);
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100000;
    regA = 32'hFFFFFFFF;
    regB = 32'h00000001; //-1+1
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100000;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b1100_0000_0000_0000_0000_0000_0000_0001; 
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100000;
    regA = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; 

    #10
    $display("\naddu");
    instruction = 32'b000000_00001_00000_00000_00000_100001;
    regA = 32'h00000001;
    regB = 32'h00000003; //3+1
    #10
    instruction = 32'b00000000001000000000000000100001;
    regA = 32'hFFFFFFFF;
    regB = 32'h00000001; 

    #10
    $display("\nand");
    instruction = 32'b000000_00001_00000_00000_00000_100100;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011; 

    #10
    $display("\nnor");
    instruction = 32'b000000_00001_00000_00000_00000_100111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011; 

    #10
    $display("\nor");
    instruction = 32'b000000_00001_00000_00000_00000_100101;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011; 

    #10
    $display("\nsll");
    instruction = 32'b000000_00000_00000_00000_00011_000000;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011;  //regA shift 3 bits left
    #10
    instruction = 32'b000000_00000_00001_00000_10000_000000;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0010_0000_0000_0000_0000_0000_0000_0011;  //regB shift 16 bits left

    #10
    $display("\nsllv");
    instruction = 32'b000000_00001_00000_00000_00011_000100;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011;  //regA << regB
    #10
    instruction = 32'b000000_00000_00001_00000_00011_000100;
    regA = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111;  //regB << regA

    #10
    $display("\nslt");
    instruction = 32'b000000_00000_00001_00000_00000_101010;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011; //rs<rt regA < regB
    #10
    instruction = 32'b000000_00001_00000_00000_00000_101010;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b1000_0000_0000_0000_0000_0000_0000_0111; //rs<rt !regB < regA

    #10
    $display("\nsltu");
    instruction = 32'b000000_00000_00001_00000_00000_101011;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0011; //rs<rt regA < regB
    #10
    instruction = 32'b000000_00001_00000_00000_00000_101011;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b1000_0000_0000_0000_0000_0000_0000_0011; //rs<rt !regB < regA

    #10
    $display("\nsra");
    instruction = 32'b000000_00000_00000_00000_00100_000011;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0010_0000_0000_0000_0000_0000_0000_0011; //regA shift 4 bits right arithmetically
    #10
    instruction = 32'b000000_00000_00001_00000_10000_000011;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0010_0000_0000_0000_0000_0000_0000_0011; //regB shift 16 bits right arithmetically

    #10
    $display("\nsrav");
    instruction = 32'b000000_00001_00000_00000_00000_000111;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0100; //regA shift 4 bits (regB) right arithmetically
    #10
    instruction = 32'b000000_00000_00001_00000_00000_000111;
    regA = 32'b1111_1111_1111_1111_1111_1111_1111_1110;
    regB = 32'b1000_0000_0000_0000_0000_0000_0000_0100; //regB shift regA bits arithmetically

    #10
    $display("\nsrl");
    instruction = 32'b000000_00000_00000_00000_00100_000010;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000; //regA shift 4 bits right logically
    #10
    instruction = 32'b000000_00000_00001_00000_00100_000010;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0100_0000_0000_0000_0000_0000_0001_1010; //regB shift 4 bits right logically

    #10
    $display("\nsrlv");
    instruction = 32'b000000_00001_00000_00000_00000_000110;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0101;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0100; //regA shift 4 bits (regB) right logically
    #10
    instruction = 32'b000000_00000_00001_00000_00000_000110;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1100; //regB shift 1 bit (regA) right logically

    #10
    $display("\nsub");
    instruction = 32'b000000_00000_00001_00000_00000_100010;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0100; //8-4
    #10
    instruction = 32'b000000_00000_00001_00000_00000_100010;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1000; //4-8
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100010;
    regA = 32'b1111_1111_1111_1111_1111_1111_1111_1000;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; //regB-regA  
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100010;
    regA = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1000_0000_0000_0000_0000_0000_0000_0000; //regB-regA  

    #10
    $display("\nsubu");
    instruction = 32'b000000_00000_00001_00000_00000_100011;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0100; //8-4 
    #10
    instruction = 32'b000000_00001_00000_00000_00000_100011;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1100_0000_0000_0000_0000_0000_0000_0000; //regB-regA    

    #10
    $display("\nxor");
    instruction = 32'b000000_00001_00000_00000_00000_100110;
    regA = 32'b0000_0000_0000_0000_0000_0000_1111_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100;

    #10
    $display("\naddi");
    instruction = 32'b001000_00000_00000_0000000000001000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; //8+8
    #10
    instruction = 32'b001000_00000_00000_1000000000000000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; 
    #10
    instruction = 32'b001000_00000_00000_1000000000000000;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; 
    #10
    instruction = 32'b001000_00001_00000_0100000000000000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0111_1111_1111_1111_1100_0000_0000_0000; //regB+immed 

    #10
    $display("\naddiu");
    instruction = 32'b001001_00000_00000_0000000000001000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; //8+8
    #10
    instruction = 32'b001001_00000_00000_1000000000000000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; 
    #10
    instruction = 32'b001001_00000_00000_1000000000000000;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_0100; 
    #10
    instruction = 32'b001001_00001_00000_0100000000000000;
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; //regB+immed 

    #10
    $display("\nandi");
    instruction = 32'b001100_00000_00000_0000000000001111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; //regA & immed

    #10
    $display("\nbeq");
    instruction = 32'b000100_00001_00000_0000000000001111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; //regA != regB flag[2]=0
    #10
    instruction = 32'b000100_00001_00000_0000000000001111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0111_1111; //regA == regB flag[2]=1

    #10
    $display("\nbne");
    instruction = 32'b000101_00001_00000_0000000000001111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0100_0000_0000_0000_0000_0000_0000_0000; //regA != regB flags[2]=0
    #10
    instruction = 32'b000101_00001_00000_0000000000001111;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0111_1111; //regA == regB flags[2]=1

    #10
    $display("\nlw");
    instruction = 32'b100011_00000_00000_0000000000000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111;  //regA+immed
    #10
    instruction = 32'b100011_00001_00000_0000000000000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111;  //regB+immed

    #10
    $display("\nori");
    instruction = 32'b001101_00000_00000_0000000010000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regA | immed
    #10
    instruction = 32'b001101_00001_00000_0000000010000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regB | immed

    #10
    $display("\nslti");
    instruction = 32'b001010_00000_00000_0000000000000001;
    regA = 32'b1000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regA < immed flags[1]=1 
    #10
    instruction = 32'b001010_00001_00000_1000000000000001;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1111_1111_1111_1111_1000_0000_0000_1111; //regB > immed flags[1]=0

    #10
    $display("\nsltiu");
    instruction = 32'b001011_00000_00000_1000000000000001;
    regA = 32'b1000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regA < immed flags[1]=1
    #10
    instruction = 32'b001011_00001_00000_0000000000000001;
    regA = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regB > immed flags[1]=0
    
    #10
    $display("\nsw");
    instruction = 32'b101011_00000_00000_0000000000000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111;  //regA+immed
    #10
    instruction = 32'b101011_00001_00000_1000000000000001;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; //regB+immed

    #10
    $display("\nxori");
    instruction = 32'b001110_00000_00000_0000000010000011;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1111; 
    #10
    instruction = 32'b001110_00001_00000_0000000010000011;
    regA = 32'b0000_0000_0000_0000_0000_0000_0111_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_1000_1111; 

end
endmodule